module main;
  initial
    begin
      $display("Happy New Year 1396!");
      $finish;
    end
endmodule
