module main;
  initial
    begin
      $display("Happy New Year 1395!");
      $finish;
    end
endmodule
